`ifndef _CONFIG_VH_
`define _CONFIG_VH_

`define cfg_divider 104  // 12 MHz / 115200 = 104.16666666666667

`endif